module rgrewallab5verilog(input [3:0]A,input [3:0]B,output reg [2:0]LED);
    reg [7:0] C;
    reg [3:0] D;
    reg [6:0] E;
    always @(A,B,C,D,E) begin
        C[0] = !A[3] && B[3];
        C[1] = A[3] && !B[3];
        C[2] = !A[2] && B[2];
        C[3] = A[2] && !B[2];
        C[4] = !A[1] && B[1];
        C[5] = A[1] && !B[1];
        C[6] = !A[0] && B[0];
        C[7] = A[0] && !B[0];

        D[0] = !(C[0] || C[1]);
        D[1] = !(C[2] || C[3]);
        D[2] = !(C[4] || C[5]);
        D[3] = !(C[6] || C[7]);

        E[0] = D[0] && C[2];
        E[1] = D[0] && C[3];
        E[2] = D[0] && D[1] && C[4];
        E[3] = D[0] && D[1] && C[5];
        E[4] = D[0] && D[1] && D[2] && C[6];
        E[5] = D[0] && D[1] && D[2] && C[7];
        E[6] = D[0] && D[1] && D[2] && D[3];

        LED[0] = C[0] || E[0] || E[2] || E[4];
        LED[1] = E[6];
        LED[2] = C[1] || E[1] || E[3] || E[5];
    end
endmodule