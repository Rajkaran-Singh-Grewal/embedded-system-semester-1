module Rgrewallab1verilog(input x,input y,output z);
assign z = x & y;
endmodule